module des_round_function
    (
        input   [31:0] R0,
        input   [47:0] K,
        output  [31:0] R1
    );

endmodule
