module des_pipeline
    (
        input clk
    );

endmodule
